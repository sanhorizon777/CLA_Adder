* C:\FOSSEE\eSim\library\SubcircuitLibrary\XOR_new\XOR_new.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 07/10/2022 18:24:41

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
SC4  Net-_SC10-Pad2_ Net-_SC3-Pad2_ GND GND sky130_fd_pr__nfet_01v8		
SC3  Net-_SC10-Pad2_ Net-_SC3-Pad2_ Net-_SC1-Pad3_ Net-_SC1-Pad3_ sky130_fd_pr__pfet_01v8		
SC2  Net-_SC1-Pad1_ Net-_SC1-Pad2_ GND GND sky130_fd_pr__nfet_01v8		
SC1  Net-_SC1-Pad1_ Net-_SC1-Pad2_ Net-_SC1-Pad3_ Net-_SC1-Pad3_ sky130_fd_pr__pfet_01v8		
U1  Net-_SC1-Pad2_ Net-_SC3-Pad2_ Net-_SC1-Pad3_ Net-_SC10-Pad1_ PORT		
SC5  Net-_SC5-Pad1_ Net-_SC3-Pad2_ Net-_SC1-Pad3_ Net-_SC1-Pad3_ sky130_fd_pr__pfet_01v8		
SC6  Net-_SC10-Pad1_ Net-_SC1-Pad1_ Net-_SC5-Pad1_ Net-_SC1-Pad3_ sky130_fd_pr__pfet_01v8		
SC9  Net-_SC10-Pad3_ Net-_SC1-Pad2_ Net-_SC1-Pad3_ Net-_SC1-Pad3_ sky130_fd_pr__pfet_01v8		
SC10  Net-_SC10-Pad1_ Net-_SC10-Pad2_ Net-_SC10-Pad3_ Net-_SC1-Pad3_ sky130_fd_pr__pfet_01v8		
SC7  Net-_SC10-Pad1_ Net-_SC1-Pad2_ Net-_SC7-Pad3_ GND sky130_fd_pr__nfet_01v8		
SC11  Net-_SC10-Pad1_ Net-_SC10-Pad2_ Net-_SC11-Pad3_ GND sky130_fd_pr__nfet_01v8		
SC8  Net-_SC7-Pad3_ Net-_SC3-Pad2_ GND GND sky130_fd_pr__nfet_01v8		
SC12  Net-_SC11-Pad3_ Net-_SC1-Pad1_ GND GND sky130_fd_pr__nfet_01v8		

.end
